magic
tech scmos
timestamp 1715137965
<< metal1 >>
rect 2541 1331 2571 1335
rect 2542 1279 2563 1283
rect 72 1113 101 1117
rect 1359 1026 1716 1030
rect 1720 1026 1721 1030
rect 1359 1018 1708 1022
rect 1712 1018 1721 1022
rect 1359 1010 1700 1014
rect 1704 1010 1721 1014
rect 1359 1002 1692 1006
rect 1696 1002 1721 1006
rect 1359 994 1684 998
rect 1688 994 1721 998
rect 1359 986 1676 990
rect 1680 986 1721 990
rect 1359 978 1668 982
rect 1672 978 1721 982
rect 1359 970 1660 974
rect 1664 970 1721 974
rect 2264 877 2571 881
rect 2238 825 2563 829
rect 10 36 14 40
rect 10 28 14 32
rect 10 20 14 24
rect 10 12 14 16
<< m2contact >>
rect 2571 1331 2575 1335
rect 2563 1279 2567 1283
rect 32 1136 36 1140
rect 1235 1123 1239 1127
rect 68 1113 72 1117
rect 101 1113 105 1117
rect 1227 1115 1231 1119
rect 1219 1107 1223 1111
rect 1211 1099 1215 1103
rect 1716 1026 1720 1030
rect 1708 1018 1712 1022
rect 1700 1010 1704 1014
rect 1692 1002 1696 1006
rect 1684 994 1688 998
rect 1676 986 1680 990
rect 1668 978 1672 982
rect 1660 970 1664 974
rect 2571 877 2575 881
rect 2563 825 2567 829
<< metal2 >>
rect 618 1185 622 1189
rect 32 868 36 1136
rect 101 1117 105 1179
rect 1211 1146 1215 1150
rect 273 1123 277 1127
rect 281 1123 285 1126
rect 289 1123 293 1126
rect 297 1122 301 1126
rect 68 868 72 1113
rect 1660 974 1664 1030
rect 1660 885 1664 970
rect 1668 982 1672 1030
rect 1668 885 1672 978
rect 1676 990 1680 1030
rect 1676 885 1680 986
rect 1684 998 1688 1030
rect 1684 885 1688 994
rect 1692 1006 1696 1030
rect 1692 885 1696 1002
rect 1700 1014 1704 1030
rect 1700 885 1704 1010
rect 1708 1022 1712 1030
rect 1708 885 1712 1018
rect 1716 885 1720 1026
rect 2563 829 2567 1279
rect 2571 881 2575 1331
rect 2605 1161 2609 1165
rect 2613 1161 2617 1165
rect 2621 1161 2625 1165
rect 2629 1161 2633 1165
rect 2637 1161 2641 1165
rect 2645 1161 2649 1165
rect 2653 1161 2657 1165
rect 2661 1161 2665 1165
rect 2266 12 2270 16
rect 2274 12 2278 16
rect 2282 12 2286 16
rect 2290 12 2294 16
rect 2298 12 2302 16
rect 2306 12 2310 16
rect 2314 12 2318 16
rect 2322 12 2326 16
use VelocityDetector  VelocityDetector_0
timestamp 1715137965
transform 1 0 9 0 1 1156
box -20 -186 2656 1091
use pvaPosition  pvaPosition_0
timestamp 1715124547
transform 1 0 0 0 1 4
box 0 -4 2326 941
<< labels >>
rlabel metal1 12 30 12 30 1 RST
rlabel metal1 12 22 12 22 1 CLK
rlabel metal1 12 14 12 14 1 B
rlabel metal1 12 38 12 38 1 A
rlabel metal2 2655 1163 2655 1163 1 V1
rlabel metal2 2647 1163 2647 1163 1 V2
rlabel metal2 2639 1163 2639 1163 1 V3
rlabel metal2 2631 1163 2631 1163 1 V4
rlabel metal2 2663 1163 2663 1163 1 V0
rlabel metal2 2623 1163 2623 1163 1 V5
rlabel metal2 2615 1163 2615 1163 1 V6
rlabel metal2 2607 1163 2607 1163 1 V7
rlabel m2contact 2565 827 2565 827 1 VSS
rlabel m2contact 2573 879 2573 879 1 VDD
rlabel metal2 2324 14 2324 14 1 P7
rlabel metal2 2316 14 2316 14 1 P6
rlabel metal2 2308 14 2308 14 1 P5
rlabel metal2 2300 14 2300 14 1 P4
rlabel metal2 2292 14 2292 14 1 P3
rlabel metal2 2284 14 2284 14 1 P2
rlabel metal2 2276 14 2276 14 1 P1
rlabel metal2 2268 14 2268 14 1 P0
rlabel metal2 299 1124 299 1124 1 C0
rlabel metal2 291 1124 291 1124 1 C1
rlabel metal2 283 1124 283 1124 1 C2
rlabel metal2 275 1125 275 1125 1 C3
rlabel m2contact 1213 1101 1213 1101 1 X0
rlabel m2contact 1221 1109 1221 1109 1 X1
rlabel m2contact 1229 1117 1229 1117 1 X2
rlabel m2contact 1237 1125 1237 1125 1 X3
rlabel metal2 620 1187 620 1187 1 NOR4
<< end >>
