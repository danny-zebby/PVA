magic
tech scmos
timestamp 1714614791
<< metal1 >>
rect -32 773 505 777
rect 509 773 533 777
rect -36 765 -28 769
rect -24 765 513 769
rect 517 765 533 769
rect -36 757 -20 761
rect -16 757 521 761
rect 525 757 533 761
rect -36 749 -12 753
rect -8 749 529 753
rect 300 668 306 672
rect 467 668 473 672
rect 477 668 533 672
rect 300 660 306 664
rect 300 576 306 580
rect 467 576 481 580
rect 485 576 533 580
rect 300 568 306 572
rect 300 484 306 488
rect 467 484 489 488
rect 493 484 533 488
rect 300 476 306 480
rect 300 392 306 396
rect 467 392 497 396
rect 501 392 533 396
rect 300 384 306 388
rect -32 356 8 360
rect 224 357 228 361
rect 300 300 306 304
rect 467 300 505 304
rect 509 300 533 304
rect 232 292 306 296
rect -24 248 8 252
rect 224 249 236 253
rect 300 208 306 212
rect 467 208 513 212
rect 517 208 533 212
rect 240 200 306 204
rect -16 140 8 144
rect 224 141 244 145
rect 300 116 306 120
rect 467 116 521 120
rect 525 116 533 120
rect 248 108 306 112
rect 221 92 288 96
rect 292 84 306 88
rect 222 40 296 44
rect -8 32 8 36
rect 224 33 252 37
rect 300 32 309 36
rect 292 24 306 28
rect 467 24 529 28
rect 256 16 306 20
rect 300 8 328 12
<< m2contact >>
rect -36 773 -32 777
rect 505 773 509 777
rect -28 765 -24 769
rect 513 765 517 769
rect -20 757 -16 761
rect 521 757 525 761
rect -12 749 -8 753
rect 529 749 533 753
rect 296 668 300 672
rect 473 668 477 672
rect 296 660 300 664
rect 296 576 300 580
rect 481 576 485 580
rect 296 568 300 572
rect 296 484 300 488
rect 489 484 493 488
rect 296 476 300 480
rect 296 392 300 396
rect 497 392 501 396
rect 296 384 300 388
rect -36 356 -32 360
rect 228 357 232 361
rect 296 300 300 304
rect 505 300 509 304
rect 228 292 232 296
rect -28 248 -24 252
rect 236 249 240 253
rect 296 208 300 212
rect 513 208 517 212
rect 236 200 240 204
rect -20 140 -16 144
rect 244 141 248 145
rect 296 116 300 120
rect 521 116 525 120
rect 244 108 248 112
rect 288 92 292 96
rect 288 84 292 88
rect 296 40 300 44
rect -12 32 -8 36
rect 252 33 256 37
rect 296 32 300 36
rect 288 24 292 28
rect 529 24 533 28
rect 252 16 256 20
rect 296 8 300 12
<< metal2 >>
rect -36 360 -32 773
rect -36 -11 -32 356
rect -28 769 -24 777
rect -28 252 -24 765
rect -28 -11 -24 248
rect -20 761 -16 777
rect -20 144 -16 757
rect -20 -11 -16 140
rect -12 753 -8 777
rect -12 36 -8 749
rect 473 672 477 777
rect 296 664 300 668
rect 296 580 300 660
rect 296 572 300 576
rect 296 488 300 568
rect 296 480 300 484
rect 296 396 300 476
rect 296 388 300 392
rect -12 -11 -8 32
rect 228 296 232 357
rect 20 0 24 4
rect 56 0 60 4
rect 228 -27 232 292
rect 296 304 300 384
rect 236 204 240 249
rect 236 -27 240 200
rect 296 212 300 300
rect 244 112 248 141
rect 244 -27 248 108
rect 296 120 300 208
rect 288 88 292 92
rect 252 20 256 33
rect 288 28 292 84
rect 296 44 300 116
rect 296 36 300 40
rect 252 -27 256 16
rect 296 12 300 32
rect 473 0 477 668
rect 481 580 485 777
rect 481 0 485 576
rect 489 488 493 777
rect 489 0 493 484
rect 497 396 501 777
rect 497 0 501 392
rect 505 304 509 773
rect 505 0 509 300
rect 513 769 517 777
rect 513 212 517 765
rect 513 0 517 208
rect 521 761 525 777
rect 521 120 525 757
rect 521 0 525 116
rect 529 753 533 777
rect 529 28 533 749
rect 529 0 533 24
use 8BitAdder  8BitAdder_0
timestamp 1714603105
transform 1 0 306 0 1 32
box -6 -32 165 706
use Reg4  Reg4_0
timestamp 1711922858
transform 1 0 0 0 1 0
box 0 0 228 432
<< labels >>
rlabel metal2 22 2 22 2 1 RST
rlabel metal2 58 2 58 2 1 CLK
rlabel metal2 254 -25 254 -25 1 Y0
rlabel metal2 246 -25 246 -25 1 Y1
rlabel metal2 238 -25 238 -25 1 Y2
rlabel metal2 230 -25 230 -25 1 Y3
rlabel m2contact 298 34 298 34 1 VSS
rlabel metal2 290 34 290 34 1 VDD
<< end >>
