magic
tech scmos
timestamp 1714623832
<< metal1 >>
rect 240 988 696 992
rect 700 988 728 992
rect 232 980 704 984
rect 708 980 728 984
rect 324 960 328 961
rect 222 956 236 960
rect 240 956 328 960
rect 222 904 228 908
rect 232 904 322 908
rect 317 897 324 901
rect -74 788 8 792
rect 224 789 252 793
rect 256 789 324 793
rect 540 790 552 794
rect 556 790 612 794
rect 700 787 718 791
rect 696 735 704 739
rect 708 735 718 739
rect -78 680 -70 684
rect -66 680 8 684
rect 224 681 260 685
rect 264 681 324 685
rect 540 682 560 686
rect 564 682 612 686
rect -78 572 -62 576
rect -58 572 8 576
rect 224 573 268 577
rect 272 573 324 577
rect 540 574 568 578
rect 572 574 612 578
rect -78 464 -54 468
rect -50 464 8 468
rect 224 465 276 469
rect 280 465 324 469
rect 540 466 576 470
rect 580 466 612 470
rect -78 356 -46 360
rect -42 356 8 360
rect 224 357 284 361
rect 288 357 324 361
rect 540 358 584 362
rect 588 358 612 362
rect -78 248 -38 252
rect -34 248 8 252
rect 224 249 292 253
rect 296 249 324 253
rect 540 250 592 254
rect 596 250 612 254
rect 636 185 718 189
rect -78 140 -30 144
rect -26 140 8 144
rect 224 141 300 145
rect 304 141 324 145
rect 540 142 600 146
rect 604 142 612 146
rect 556 90 648 94
rect 564 82 656 86
rect 572 74 664 78
rect 580 66 672 70
rect 588 58 680 62
rect 596 50 688 54
rect 604 42 696 46
rect -78 32 -22 36
rect -18 32 8 36
rect 224 33 308 37
rect 312 33 324 37
rect 540 34 608 38
rect 612 34 704 38
rect 28 -20 56 -16
rect 60 -20 372 -16
rect 24 -28 336 -24
rect 249 -41 252 -37
rect 256 -41 967 -37
rect 971 -41 1027 -37
rect 249 -49 260 -45
rect 264 -49 975 -45
rect 979 -49 1027 -45
rect 249 -57 268 -53
rect 272 -57 983 -53
rect 987 -57 1027 -53
rect 249 -65 276 -61
rect 280 -65 991 -61
rect 995 -65 1027 -61
rect 249 -73 284 -69
rect 288 -73 999 -69
rect 1003 -73 1027 -69
rect 249 -81 292 -77
rect 296 -81 1007 -77
rect 1011 -81 1027 -77
rect 249 -89 300 -85
rect 304 -89 1015 -85
rect 1019 -89 1027 -85
rect 249 -97 308 -93
rect 312 -97 1023 -93
<< m2contact >>
rect 236 988 240 992
rect 696 988 700 992
rect 228 980 232 984
rect 704 980 708 984
rect 236 956 240 960
rect 228 904 232 908
rect -78 788 -74 792
rect 252 789 256 793
rect 552 790 556 794
rect 696 787 700 791
rect 704 735 708 739
rect -70 680 -66 684
rect 260 681 264 685
rect 560 682 564 686
rect -62 572 -58 576
rect 268 573 272 577
rect 568 574 572 578
rect -54 464 -50 468
rect 276 465 280 469
rect 576 466 580 470
rect -46 356 -42 360
rect 284 357 288 361
rect 584 358 588 362
rect -38 248 -34 252
rect 292 249 296 253
rect 592 250 596 254
rect 632 185 636 189
rect -30 140 -26 144
rect 300 141 304 145
rect 600 142 604 146
rect 552 90 556 94
rect 648 90 652 94
rect 560 82 564 86
rect 656 82 660 86
rect 568 74 572 78
rect 664 74 668 78
rect 576 66 580 70
rect 672 66 676 70
rect 584 58 588 62
rect 680 58 684 62
rect 592 50 596 54
rect 688 50 692 54
rect 600 42 604 46
rect 696 42 700 46
rect -22 32 -18 36
rect 308 33 312 37
rect 608 34 612 38
rect 704 34 708 38
rect 56 -20 60 -16
rect 372 -20 376 -16
rect 20 -28 24 -24
rect 336 -28 340 -24
rect 252 -41 256 -37
rect 967 -41 971 -37
rect 260 -49 264 -45
rect 975 -49 979 -45
rect 268 -57 272 -53
rect 983 -57 987 -53
rect 276 -65 280 -61
rect 991 -65 995 -61
rect 284 -73 288 -69
rect 999 -73 1003 -69
rect 292 -81 296 -77
rect 1007 -81 1011 -77
rect 300 -89 304 -85
rect 1015 -89 1019 -85
rect 308 -97 312 -93
rect 1023 -97 1027 -93
<< metal2 >>
rect 228 908 232 980
rect 236 960 240 988
rect 252 793 256 960
rect -78 -46 -74 788
rect -70 684 -66 792
rect -70 -46 -66 680
rect -62 576 -58 792
rect -62 -46 -58 572
rect -54 468 -50 792
rect -54 -46 -50 464
rect -46 360 -42 792
rect -46 -46 -42 356
rect -38 252 -34 792
rect -38 -46 -34 248
rect -30 144 -26 792
rect -30 -46 -26 140
rect -22 36 -18 792
rect -22 -46 -18 32
rect 20 -24 24 0
rect 56 -16 60 1
rect 252 -37 256 789
rect 252 -99 256 -41
rect 260 685 264 960
rect 260 -45 264 681
rect 260 -99 264 -49
rect 268 577 272 960
rect 268 -53 272 573
rect 268 -99 272 -57
rect 276 469 280 960
rect 276 -61 280 465
rect 276 -99 280 -65
rect 284 361 288 960
rect 284 -69 288 357
rect 284 -99 288 -73
rect 292 253 296 960
rect 292 -77 296 249
rect 292 -99 296 -81
rect 300 145 304 960
rect 300 -85 304 141
rect 300 -99 304 -89
rect 308 37 312 960
rect 552 94 556 790
rect 560 686 564 794
rect 560 86 564 682
rect 568 578 572 794
rect 568 78 572 574
rect 576 470 580 794
rect 576 70 580 466
rect 584 362 588 794
rect 584 62 588 358
rect 592 254 596 794
rect 592 54 596 250
rect 600 146 604 794
rect 600 46 604 142
rect 608 38 612 794
rect 696 791 700 988
rect 704 739 708 980
rect 664 78 668 85
rect 672 70 676 85
rect 680 62 684 85
rect 688 54 692 85
rect 696 46 700 85
rect 704 38 708 85
rect 308 -93 312 33
rect 336 -24 340 4
rect 372 -16 376 7
rect 967 -37 971 6
rect 967 -97 971 -41
rect 975 -45 979 6
rect 975 -97 979 -49
rect 983 -53 987 6
rect 983 -97 987 -57
rect 991 -61 995 6
rect 991 -97 995 -65
rect 999 -69 1003 6
rect 999 -97 1003 -73
rect 1007 -77 1011 6
rect 1007 -97 1011 -81
rect 1015 -85 1019 6
rect 1015 -97 1019 -89
rect 1023 -93 1027 6
rect 1228 -39 1232 75
rect 1236 -39 1240 75
rect 1244 -39 1248 75
rect 1252 -39 1256 75
rect 1260 -39 1264 75
rect 1268 -39 1272 75
rect 1276 -39 1280 75
rect 1284 -39 1288 75
rect 308 -99 312 -97
use Reg8  Reg8_0
timestamp 1711923903
transform 1 0 0 0 1 0
box 0 0 228 972
use Reg8  Reg8_1
timestamp 1711923903
transform 1 0 316 0 1 1
box 0 0 228 972
use SUB8  SUB8_0
timestamp 1714615921
transform 1 0 1045 0 1 109
box -413 -109 243 738
<< labels >>
rlabel m2contact 22 -26 22 -26 1 RST
rlabel metal1 30 -18 30 -18 1 EN
rlabel metal2 1286 -37 1286 -37 1 Y0
rlabel metal2 1278 -37 1278 -37 1 Y1
rlabel metal2 1270 -37 1270 -37 1 Y2
rlabel metal2 1262 -37 1262 -37 1 Y3
rlabel metal2 1254 -37 1254 -37 1 Y4
rlabel metal2 1246 -37 1246 -37 1 Y5
rlabel metal2 1238 -37 1238 -37 1 Y6
rlabel metal2 1230 -37 1230 -37 1 Y7
rlabel metal2 -28 -44 -28 -44 1 A1
rlabel metal2 -20 -44 -20 -44 1 A0
rlabel metal2 -36 -44 -36 -44 1 A2
rlabel metal2 -44 -44 -44 -44 1 A3
rlabel metal2 -52 -44 -52 -44 1 A4
rlabel metal2 -60 -44 -60 -44 1 A5
rlabel metal2 -68 -44 -68 -44 1 A6
rlabel metal2 -76 -44 -76 -44 1 A7
rlabel metal1 235 958 235 958 1 VDD
rlabel metal1 234 906 234 906 1 VSS
rlabel metal1 250 -95 250 -95 1 X0
rlabel metal1 250 -87 250 -87 1 X1
rlabel metal1 250 -79 250 -79 1 X2
rlabel metal1 250 -71 250 -71 1 X3
rlabel metal1 250 -63 250 -63 1 X4
rlabel metal1 250 -55 250 -55 1 X5
rlabel metal1 250 -47 250 -47 1 X6
rlabel metal1 250 -39 250 -39 1 X7
<< end >>
