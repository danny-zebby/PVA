magic
tech scmos
timestamp 1711564571
<< nwell >>
rect -6 38 46 62
<< ntransistor >>
rect 7 8 9 12
rect 15 8 17 12
rect 23 8 25 12
rect 31 8 33 12
<< ptransistor >>
rect 7 44 9 48
rect 15 44 17 48
rect 23 44 25 48
rect 31 44 33 48
<< ndiffusion >>
rect 6 8 7 12
rect 9 8 10 12
rect 14 8 15 12
rect 17 8 18 12
rect 22 8 23 12
rect 25 8 26 12
rect 30 8 31 12
rect 33 8 34 12
<< pdiffusion >>
rect 6 44 7 48
rect 9 44 15 48
rect 17 44 23 48
rect 25 44 31 48
rect 33 44 34 48
<< ndcontact >>
rect 2 8 6 12
rect 10 8 14 12
rect 18 8 22 12
rect 26 8 30 12
rect 34 8 38 12
<< pdcontact >>
rect 2 44 6 48
rect 34 44 38 48
<< psubstratepcontact >>
rect 2 0 6 4
<< nsubstratencontact >>
rect 2 52 6 56
<< polysilicon >>
rect 7 48 9 50
rect 15 48 17 50
rect 23 48 25 50
rect 31 48 33 50
rect 7 28 9 44
rect 15 28 17 44
rect 23 28 25 44
rect 31 28 33 44
rect 7 12 9 24
rect 15 12 17 24
rect 23 12 25 24
rect 31 12 33 24
rect 7 6 9 8
rect 15 6 17 8
rect 23 6 25 8
rect 31 6 33 8
<< polycontact >>
rect 6 24 10 28
rect 14 24 18 28
rect 22 24 26 28
rect 30 24 34 28
<< metal1 >>
rect 0 52 2 56
rect 6 52 40 56
rect 2 48 6 52
rect 34 40 38 44
rect 2 16 34 20
rect 2 12 6 16
rect 18 12 22 16
rect 34 12 38 16
rect 10 4 14 8
rect 26 4 30 8
rect 0 0 2 4
rect 6 0 40 4
<< m2contact >>
rect 34 36 38 40
rect 34 16 38 20
<< metal2 >>
rect 34 20 38 36
<< labels >>
rlabel psubstratepcontact 4 2 4 2 1 VSS
rlabel nsubstratencontact 4 54 4 54 1 VDD
rlabel polycontact 8 26 8 26 1 A
rlabel polycontact 16 26 16 26 1 B
rlabel polycontact 24 26 24 26 1 C
rlabel polycontact 32 26 32 26 1 D
rlabel m2contact 36 18 36 18 1 Y
<< end >>
