magic
tech scmos
timestamp 1714882249
<< metal1 >>
rect 2193 934 5410 938
rect 2193 926 5410 930
rect 2193 918 5410 922
rect 2193 910 5410 914
rect 2193 902 5410 906
rect 2193 894 5410 898
rect 2193 886 5410 890
rect 2193 878 5410 882
rect 952 343 997 347
rect 960 214 987 218
rect -60 72 18 76
rect -60 64 18 68
rect -60 56 18 60
rect 977 58 992 62
rect -60 48 18 52
rect 977 28 981 58
rect 920 24 981 28
rect 986 20 990 54
rect 928 16 990 20
rect 2639 15 2843 19
rect 2639 1 2643 15
rect 2654 7 5410 11
rect 2025 -3 2643 1
rect 2650 -1 2658 3
rect 2662 -1 5410 3
rect 4 -11 2189 -7
rect 2670 -9 5410 -5
rect -4 -19 2197 -15
rect 2678 -17 5410 -13
rect -12 -27 2205 -23
rect 2686 -25 5410 -21
rect -20 -35 2213 -31
rect 2694 -33 5410 -29
rect -28 -43 2221 -39
rect 2702 -41 5410 -37
rect -36 -51 2229 -47
rect 2710 -49 5410 -45
rect -44 -59 2237 -55
rect -52 -67 2245 -63
rect 5351 -882 5410 -878
rect 5359 -890 5410 -886
rect 5367 -898 5410 -894
rect 5375 -906 5410 -902
rect 5383 -914 5410 -910
rect 5391 -922 5410 -918
rect 5399 -930 5410 -926
rect 5399 -938 5410 -934
rect 24 -1192 52 -1188
rect 1657 -1192 2752 -1189
rect -52 -1302 34 -1298
rect 2654 -1300 2740 -1296
rect -44 -1310 41 -1306
rect 2662 -1308 2749 -1304
rect -36 -1318 48 -1314
rect 2670 -1316 2756 -1312
rect -28 -1326 56 -1322
rect 2678 -1324 2765 -1320
rect -20 -1334 64 -1330
rect 2686 -1332 2772 -1328
rect -12 -1342 71 -1338
rect 2694 -1340 2780 -1336
rect -4 -1350 37 -1346
rect 2702 -1348 2789 -1344
rect 4 -1358 35 -1354
rect 2710 -1356 2796 -1352
<< m2contact >>
rect 948 343 952 347
rect 956 214 960 218
rect 575 168 579 172
rect 146 56 150 60
rect 2843 15 2847 19
rect 2650 7 2654 11
rect 2658 -1 2662 3
rect 0 -11 4 -7
rect 2189 -11 2193 -7
rect 2666 -9 2670 -5
rect -8 -19 -4 -15
rect 2197 -19 2201 -15
rect 2674 -17 2678 -13
rect -16 -27 -12 -23
rect 2205 -27 2209 -23
rect 2682 -25 2686 -21
rect -24 -35 -20 -31
rect 2213 -35 2217 -31
rect 2690 -33 2694 -29
rect -32 -43 -28 -39
rect 2221 -43 2225 -39
rect 2698 -41 2702 -37
rect -40 -51 -36 -47
rect 2229 -51 2233 -47
rect 2706 -49 2710 -45
rect -48 -59 -44 -55
rect 2237 -59 2241 -55
rect -56 -67 -52 -63
rect 2245 -67 2249 -63
rect 1430 -113 1434 -109
rect 4239 -115 4243 -111
rect 5347 -882 5351 -878
rect 3412 -887 3416 -883
rect 5355 -890 5359 -886
rect 5363 -898 5367 -894
rect 5371 -906 5375 -902
rect 5379 -914 5383 -910
rect 5387 -922 5391 -918
rect 5395 -930 5399 -926
rect 713 -997 717 -993
rect 20 -1192 24 -1188
rect -56 -1302 -52 -1298
rect 2650 -1300 2654 -1296
rect -48 -1310 -44 -1306
rect 2658 -1308 2662 -1304
rect -40 -1318 -36 -1314
rect 2666 -1316 2670 -1312
rect -32 -1326 -28 -1322
rect 2674 -1324 2678 -1320
rect -24 -1334 -20 -1330
rect 2682 -1332 2686 -1328
rect -16 -1342 -12 -1338
rect 2690 -1340 2694 -1336
rect -8 -1350 -4 -1346
rect 2698 -1348 2702 -1344
rect 0 -1358 4 -1354
rect 2706 -1356 2710 -1352
<< metal2 >>
rect 948 188 952 343
rect -56 -1298 -52 -67
rect -48 -1306 -44 -59
rect -40 -1314 -36 -51
rect -32 -1322 -28 -43
rect -24 -1330 -20 -35
rect -16 -1338 -12 -27
rect -8 -1346 -4 -19
rect 0 -1354 4 -11
rect 20 -1188 24 28
rect 146 -713 150 56
rect 2189 -7 2193 13
rect 2197 -15 2201 13
rect 2205 -23 2209 13
rect 2213 -31 2217 13
rect 2221 -39 2225 13
rect 2229 -47 2233 13
rect 2237 -55 2241 13
rect 2245 -63 2249 13
rect 2650 -1296 2654 7
rect 2658 -1304 2662 -1
rect 2666 -1312 2670 -9
rect 2674 -1320 2678 -17
rect 2682 -1328 2686 -25
rect 2690 -1336 2694 -33
rect 2690 -1356 2694 -1340
rect 2698 -1344 2702 -41
rect 2698 -1356 2702 -1348
rect 2706 -1352 2710 -49
rect 2843 -711 2847 15
rect 2843 -715 2846 -711
<< m3contact >>
rect 587 888 591 892
rect 2105 870 2109 874
rect 152 848 156 852
rect 579 168 583 172
rect 2161 169 2165 173
rect 1430 -109 1434 -105
rect 709 -997 713 -993
rect 4243 -115 4247 -111
rect 3408 -887 3412 -883
<< metal3 >>
rect 1323 939 1463 940
rect 2252 939 5410 940
rect -55 933 5410 939
rect -60 892 5410 933
rect -60 888 587 892
rect 591 888 5410 892
rect -60 874 5410 888
rect -60 870 2105 874
rect 2109 870 5410 874
rect -60 852 5410 870
rect -60 848 152 852
rect 156 848 5410 852
rect -60 814 5410 848
rect -60 811 2253 814
rect -60 -792 80 811
rect 578 172 718 706
rect 578 168 579 172
rect 583 168 718 172
rect 578 -876 718 168
rect 1323 -105 1463 811
rect 1323 -109 1430 -105
rect 1434 -109 1463 -105
rect 1323 -785 1463 -109
rect 2106 173 2246 706
rect 2106 169 2161 173
rect 2165 169 2246 173
rect 2106 -876 2246 169
rect 3023 -876 3427 456
rect 4125 -111 4867 814
rect 4125 -115 4243 -111
rect 4247 -115 4867 -111
rect 4125 -815 4867 -115
rect 5107 -876 5410 653
rect -67 -883 5410 -876
rect -67 -887 3408 -883
rect 3412 -887 5410 -883
rect -67 -993 5410 -887
rect -67 -997 709 -993
rect 713 -997 5410 -993
rect -67 -1359 5410 -997
use PositionPart  PositionPart_0
timestamp 1714633149
transform 1 0 1064 0 1 114
box -81 -117 1185 824
use VelocityDetector  VelocityDetector_0
timestamp 1714633149
transform 1 0 54 0 1 -1172
box -20 -186 2656 1091
use VelocityDetector  VelocityDetector_1
timestamp 1714633149
transform 1 0 2751 0 1 -1170
box -20 -186 2656 1091
use directionDetector  directionDetector_0
timestamp 1712454563
transform 1 0 0 0 1 48
box 0 -48 960 856
<< labels >>
rlabel metal2 2652 -1161 2652 -1161 7 Y0
rlabel metal2 2652 -1110 2652 -1110 1 Y0
rlabel metal2 2652 -996 2652 -996 7 Y0
rlabel metal2 2660 -1161 2660 -1161 7 Y0
rlabel metal2 2660 -1110 2660 -1110 1 Y0
rlabel metal2 2660 -996 2660 -996 7 Y0
rlabel metal2 2660 -1161 2660 -1161 1 Y7
rlabel metal2 2660 -1110 2660 -1110 1 Y7
rlabel metal2 2660 -996 2660 -996 1 Y7
rlabel metal2 2668 -1161 2668 -1161 7 Y0
rlabel metal2 2668 -1110 2668 -1110 1 Y0
rlabel metal2 2668 -996 2668 -996 7 Y0
rlabel metal2 2668 -1161 2668 -1161 1 Y7
rlabel metal2 2668 -1110 2668 -1110 1 Y7
rlabel metal2 2668 -996 2668 -996 1 Y7
rlabel metal2 2676 -1161 2676 -1161 7 Y0
rlabel metal2 2676 -1110 2676 -1110 1 Y0
rlabel metal2 2676 -996 2676 -996 7 Y0
rlabel metal2 2676 -1161 2676 -1161 1 Y7
rlabel metal2 2676 -1110 2676 -1110 1 Y7
rlabel metal2 2676 -996 2676 -996 1 Y7
rlabel metal2 2684 -1161 2684 -1161 7 Y0
rlabel metal2 2684 -1110 2684 -1110 1 Y0
rlabel metal2 2684 -996 2684 -996 7 Y0
rlabel metal2 2684 -1161 2684 -1161 1 Y7
rlabel metal2 2684 -1110 2684 -1110 1 Y7
rlabel metal2 2684 -996 2684 -996 1 Y7
rlabel metal2 2692 -1161 2692 -1161 7 Y0
rlabel metal2 2692 -1110 2692 -1110 1 Y0
rlabel metal2 2692 -996 2692 -996 7 Y0
rlabel metal2 2692 -1161 2692 -1161 1 Y7
rlabel metal2 2692 -1110 2692 -1110 1 Y7
rlabel metal2 2692 -996 2692 -996 1 Y7
rlabel metal2 2700 -1161 2700 -1161 7 Y0
rlabel metal2 2700 -1110 2700 -1110 1 Y0
rlabel metal2 2700 -996 2700 -996 7 Y0
rlabel metal2 2700 -1161 2700 -1161 1 Y7
rlabel metal2 2700 -1110 2700 -1110 1 Y7
rlabel metal2 2700 -996 2700 -996 1 Y7
rlabel metal2 2708 -1161 2708 -1161 7 Y0
rlabel metal2 2708 -1110 2708 -1110 1 Y0
rlabel metal2 2708 -996 2708 -996 7 Y0
rlabel metal2 2708 -1161 2708 -1161 1 Y7
rlabel metal2 2708 -1110 2708 -1110 1 Y7
rlabel metal2 2708 -996 2708 -996 1 Y7
rlabel metal3 3231 217 3231 217 1 VSS
rlabel metal3 4370 174 4370 174 1 VDD
rlabel metal1 -59 74 -59 74 1 A
rlabel metal1 -59 66 -59 66 1 RST
rlabel metal1 -59 58 -59 58 1 CLK
rlabel metal1 -59 50 -59 50 1 B
rlabel metal1 5409 936 5409 936 6 P7
rlabel metal1 5409 928 5409 928 7 P6
rlabel metal1 5409 920 5409 920 7 P5
rlabel metal1 5409 912 5409 912 7 P4
rlabel metal1 5409 904 5409 904 7 P3
rlabel metal1 5409 896 5409 896 7 P2
rlabel metal1 5409 888 5409 888 7 P1
rlabel metal1 5409 880 5409 880 7 P0
rlabel metal1 5409 9 5409 9 7 V7
rlabel metal1 5409 1 5409 1 7 V6
rlabel metal1 5409 -7 5409 -7 7 V5
rlabel metal1 5409 -15 5409 -15 7 V4
rlabel metal1 5409 -23 5409 -23 7 V3
rlabel metal1 5409 -31 5409 -31 7 V2
rlabel metal1 5409 -39 5409 -39 7 V1
rlabel metal1 5409 -47 5409 -47 7 V0
rlabel metal1 5409 -936 5409 -936 7 A0
rlabel metal1 5409 -928 5409 -928 7 A1
rlabel metal1 5409 -920 5409 -920 7 A2
rlabel metal1 5409 -912 5409 -912 7 A3
rlabel metal1 5409 -904 5409 -904 7 A4
rlabel metal1 5409 -896 5409 -896 7 A5
rlabel metal1 5409 -888 5409 -888 7 A6
rlabel metal1 5409 -880 5409 -880 7 A7
<< end >>
