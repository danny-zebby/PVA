magic
tech scmos
timestamp 1714615249
use DFFMUX  DFFMUX_0
timestamp 1714612951
transform 1 0 0 0 1 0
box -4 -48 366 68
use DFFMUX  DFFMUX_1
timestamp 1714612951
transform 1 0 0 0 1 108
box -4 -48 366 68
use DFFMUX  DFFMUX_2
timestamp 1714612951
transform 1 0 0 0 1 216
box -4 -48 366 68
use DFFMUX  DFFMUX_3
timestamp 1714612951
transform 1 0 0 0 1 325
box -4 -48 366 68
use DFFMUX  DFFMUX_4
timestamp 1714612951
transform 1 0 0 0 1 433
box -4 -48 366 68
use DFFMUX  DFFMUX_5
timestamp 1714612951
transform 1 0 0 0 1 541
box -4 -48 366 68
use DFFMUX  DFFMUX_6
timestamp 1714612951
transform 1 0 0 0 1 649
box -4 -48 366 68
use DFFMUX  DFFMUX_7
timestamp 1714612951
transform 1 0 0 0 1 757
box -4 -48 366 68
<< labels >>
rlabel metal1 1 -22 1 -22 3 D0
rlabel metal1 1 -6 1 -6 3 en
rlabel metal1 1 2 1 2 3 VSS
rlabel metal1 1 54 1 54 3 VDD
rlabel metal1 1 86 1 86 3 D1
rlabel metal1 1 194 1 194 3 D2
rlabel metal1 1 303 1 303 3 D3
rlabel metal1 1 411 1 411 3 D4
rlabel metal1 1 519 1 519 3 D5
rlabel metal1 1 627 1 627 3 D6
rlabel metal1 1 735 1 735 3 D7
rlabel metal1 151 -14 151 -14 1 RST
rlabel metal1 151 -22 151 -22 1 CLK
rlabel metal1 359 751 359 751 1 Q7
rlabel metal1 359 742 359 742 1 Q7b
rlabel metal1 359 643 359 643 1 Q6
rlabel metal1 359 634 359 634 1 Q6b
rlabel metal1 359 535 359 535 1 Q5
rlabel metal1 359 526 359 526 1 Q5b
rlabel metal1 359 427 359 427 1 Q4
rlabel metal1 359 418 359 418 1 Q4b
rlabel metal1 359 319 359 319 1 Q3
rlabel metal1 359 310 359 310 1 Q3b
rlabel metal1 359 210 359 210 1 Q2
rlabel metal1 359 201 359 201 1 Q2b
rlabel metal1 359 102 359 102 1 Q1
rlabel metal1 359 93 359 93 1 Q1b
rlabel metal1 359 -6 359 -6 1 Q0
rlabel metal1 359 -15 359 -15 1 Q0b
<< end >>
