magic
tech scmos
timestamp 1711594718
<< nwell >>
rect 8 52 12 56
<< psubstratepcontact >>
rect 8 0 12 4
<< nsubstratencontact >>
rect 8 52 12 56
<< polycontact >>
rect 12 24 16 28
rect 20 24 24 28
rect 28 24 32 28
<< metal1 >>
rect 36 20 48 24
rect 52 16 56 20
use INV  INV_0
timestamp 1711561836
transform 1 0 42 0 1 0
box -4 0 20 59
use NAND3  NAND3_0
timestamp 1711593430
transform 1 0 6 0 1 0
box -6 0 42 62
<< labels >>
rlabel nsubstratencontact 10 54 10 54 1 VDD
rlabel psubstratepcontact 10 2 10 2 1 VSS
rlabel metal1 54 18 54 18 1 Y
rlabel polycontact 14 26 14 26 1 A
rlabel polycontact 22 26 22 26 1 B
rlabel polycontact 30 26 30 26 1 C
<< end >>
