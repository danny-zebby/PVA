magic
tech scmos
timestamp 1714606253
<< nwell >>
rect -213 592 -205 596
rect -213 506 -205 510
rect -213 420 -205 424
rect -213 334 -205 338
rect -213 248 -205 252
rect -213 162 -205 166
rect -213 76 -205 80
<< metal1 >>
rect -213 678 -201 682
rect -74 668 32 672
rect 149 668 183 672
rect 0 660 7 664
rect -217 642 -164 646
rect -160 642 -4 646
rect -222 626 -209 630
rect -393 618 -266 622
rect -409 610 -298 614
rect -213 592 -201 596
rect -66 576 32 580
rect 149 576 191 580
rect 2 560 7 572
rect -217 556 -156 560
rect -152 556 7 560
rect -222 540 -209 544
rect -385 532 -266 536
rect -409 524 -298 528
rect -213 506 -201 510
rect -58 484 32 488
rect 149 484 199 488
rect 2 474 6 480
rect -217 470 -148 474
rect -144 470 6 474
rect -222 454 -209 458
rect -377 446 -266 450
rect -409 438 -298 442
rect -213 420 -201 424
rect -50 392 32 396
rect 149 392 207 396
rect -217 384 -140 388
rect -136 384 9 388
rect -222 368 -209 372
rect -369 360 -266 364
rect -409 352 -298 356
rect -213 334 -201 338
rect -217 298 -132 302
rect -128 298 -104 302
rect -42 300 32 304
rect 149 300 215 304
rect 1 292 7 296
rect -128 288 6 292
rect -222 282 -209 286
rect -361 274 -298 278
rect -409 266 -298 270
rect -213 248 -201 252
rect -217 212 -124 216
rect -120 212 -104 216
rect -34 208 32 212
rect 149 208 223 212
rect -120 200 40 204
rect -222 196 -209 200
rect -353 188 -325 192
rect -409 180 -298 184
rect -213 162 -201 166
rect -217 126 -116 130
rect -112 126 -104 130
rect -26 116 19 120
rect 149 116 231 120
rect -222 110 -209 114
rect -112 108 6 112
rect -345 102 -325 106
rect -409 94 -298 98
rect -197 84 6 88
rect -213 76 -201 80
rect -217 40 -108 44
rect -205 32 6 36
rect -219 24 -209 28
rect -18 24 9 28
rect 167 24 239 28
rect -337 16 -321 20
rect -104 16 6 20
rect -409 8 -298 12
rect -197 -33 4 -29
rect 118 -69 125 -65
rect -205 -85 4 -81
rect -409 -93 47 -89
<< m2contact >>
rect -201 678 -197 682
rect -78 668 -74 672
rect 183 668 187 672
rect -4 660 0 664
rect -164 642 -160 646
rect -4 642 0 646
rect -209 626 -205 630
rect -397 618 -393 622
rect -413 610 -409 614
rect -201 592 -197 596
rect -70 576 -66 580
rect 191 576 195 580
rect -156 556 -152 560
rect -209 540 -205 544
rect -389 532 -385 536
rect -413 524 -409 528
rect -201 506 -197 510
rect -62 484 -58 488
rect 199 484 203 488
rect -148 470 -144 474
rect -209 454 -205 458
rect -381 446 -377 450
rect -413 438 -409 442
rect -201 420 -197 424
rect -54 392 -50 396
rect 207 392 211 396
rect -140 384 -136 388
rect -209 368 -205 372
rect -373 360 -369 364
rect -413 352 -409 356
rect -201 334 -197 338
rect -132 298 -128 302
rect -46 300 -42 304
rect 215 300 219 304
rect -132 288 -128 292
rect -209 282 -205 286
rect -365 274 -361 278
rect -413 266 -409 270
rect -201 248 -197 252
rect -124 212 -120 216
rect -38 208 -34 212
rect 223 208 227 212
rect -124 200 -120 204
rect -209 196 -205 200
rect -357 188 -353 192
rect -413 180 -409 184
rect -201 162 -197 166
rect -116 126 -112 130
rect -30 116 -26 120
rect 231 116 235 120
rect -209 110 -205 114
rect -116 108 -112 112
rect -349 102 -345 106
rect -413 94 -409 98
rect -201 84 -197 88
rect -201 76 -197 80
rect -108 40 -104 44
rect -209 32 -205 36
rect -209 24 -205 28
rect -22 24 -18 28
rect 239 24 243 28
rect -341 16 -337 20
rect -108 16 -104 20
rect -413 8 -409 12
rect -201 -33 -197 -29
rect 114 -69 118 -65
rect 125 -69 129 -65
rect -209 -85 -205 -81
rect 33 -85 37 -81
rect -413 -93 -409 -89
<< metal2 >>
rect -413 614 -409 619
rect -413 528 -409 610
rect -413 442 -409 524
rect -413 356 -409 438
rect -413 270 -409 352
rect -413 184 -409 266
rect -413 98 -409 180
rect -413 12 -409 94
rect -413 -89 -409 8
rect -397 -24 -393 618
rect -389 536 -385 622
rect -389 -24 -385 532
rect -381 450 -377 622
rect -381 -24 -377 446
rect -373 364 -369 622
rect -373 -24 -369 360
rect -365 278 -361 622
rect -365 -24 -361 274
rect -357 192 -353 622
rect -357 -24 -353 188
rect -349 106 -345 622
rect -349 -24 -345 102
rect -341 20 -337 622
rect -341 -24 -337 16
rect -209 544 -205 626
rect -209 458 -205 540
rect -209 372 -205 454
rect -209 286 -205 368
rect -209 200 -205 282
rect -209 114 -205 196
rect -209 36 -205 110
rect -209 28 -205 32
rect -209 -81 -205 24
rect -201 596 -197 678
rect -201 510 -197 592
rect -201 424 -197 506
rect -201 338 -197 420
rect -201 252 -197 334
rect -201 166 -197 248
rect -201 88 -197 162
rect -201 80 -197 84
rect -201 -29 -197 76
rect -164 40 -160 642
rect -156 560 -152 646
rect -156 40 -152 556
rect -148 474 -144 646
rect -148 40 -144 470
rect -140 388 -136 646
rect -140 40 -136 384
rect -132 302 -128 646
rect -132 292 -128 298
rect -132 40 -128 288
rect -124 216 -120 646
rect -124 204 -120 212
rect -124 40 -120 200
rect -116 130 -112 646
rect -116 112 -112 126
rect -116 40 -112 108
rect -108 44 -104 646
rect -108 20 -104 40
rect -78 -103 -74 668
rect -70 580 -66 668
rect -70 -103 -66 576
rect -62 488 -58 668
rect -62 -103 -58 484
rect -54 396 -50 668
rect -54 -103 -50 392
rect -46 304 -42 668
rect -46 -103 -42 300
rect -38 212 -34 668
rect -38 -103 -34 208
rect -30 120 -26 668
rect -30 -103 -26 116
rect -22 28 -18 668
rect -4 646 0 660
rect -22 -103 -18 24
rect 125 -65 129 48
rect 183 -34 187 668
rect 191 -34 195 576
rect 199 -34 203 484
rect 207 -34 211 392
rect 215 -34 219 300
rect 223 -34 227 208
rect 231 -34 235 116
rect 239 -34 243 24
use 8BitAdder  8BitAdder_0
timestamp 1713982514
transform 1 0 6 0 1 32
box -6 -32 165 706
use XOR2  XOR2_0
timestamp 1711599452
transform 1 0 -331 0 1 540
box 0 -24 126 62
use XOR2  XOR2_1
timestamp 1711599452
transform 1 0 -331 0 1 368
box 0 -24 126 62
use XOR2  XOR2_2
timestamp 1711599452
transform 1 0 -331 0 1 454
box 0 -24 126 62
use XOR2  XOR2_3
timestamp 1711599452
transform 1 0 -331 0 1 626
box 0 -24 126 62
use XOR2  XOR2_4
timestamp 1711599452
transform 1 0 -331 0 1 282
box 0 -24 126 62
use XOR2  XOR2_5
timestamp 1711599452
transform 1 0 -331 0 1 196
box 0 -24 126 62
use XOR2  XOR2_6
timestamp 1711599452
transform 1 0 -331 0 1 110
box 0 -24 126 62
use XOR2  XOR2_7
timestamp 1711599452
transform 1 0 0 0 1 -85
box 0 -24 126 62
use XOR2  XOR2_8
timestamp 1711599452
transform 1 0 -331 0 1 24
box 0 -24 126 62
<< labels >>
rlabel metal2 241 -32 241 -32 7 Y0
rlabel metal2 233 -32 233 -32 1 Y1
rlabel metal2 225 -32 225 -32 1 Y2
rlabel metal2 217 -32 217 -32 1 Y3
rlabel metal2 209 -32 209 -32 1 Y4
rlabel metal2 201 -32 201 -32 1 Y5
rlabel metal2 193 -32 193 -32 1 Y6
rlabel metal2 185 -32 185 -32 1 Y7
rlabel metal2 -20 -101 -20 -101 1 A0
rlabel metal2 -28 -101 -28 -101 1 A1
rlabel metal2 -36 -101 -36 -101 1 A2
rlabel metal2 -44 -101 -44 -101 1 A3
rlabel metal2 -52 -101 -52 -101 1 A4
rlabel metal2 -60 -101 -60 -101 1 A5
rlabel metal2 -68 -101 -68 -101 1 A6
rlabel m2contact -199 78 -199 78 1 VDD
rlabel m2contact -207 26 -207 26 1 VSS
rlabel metal2 -339 -22 -339 -22 1 B0
rlabel metal2 -347 -22 -347 -22 1 B1
rlabel metal2 -355 -22 -355 -22 1 B2
rlabel metal2 -363 -22 -363 -22 1 B3
rlabel metal2 -371 -22 -371 -22 1 B4
rlabel metal2 -379 -22 -379 -22 1 B5
rlabel metal2 -387 -22 -387 -22 1 B6
rlabel metal2 -395 -22 -395 -22 1 B7
rlabel metal2 -411 -21 -411 -21 3 SEL
rlabel metal2 -76 -101 -76 -101 1 A7
rlabel metal1 -215 130 -215 130 1 Y
rlabel metal1 -215 216 -215 216 1 Y
rlabel metal1 -215 302 -215 302 1 Y
rlabel metal1 -215 388 -215 388 1 Y
rlabel metal1 -215 474 -215 474 1 Y
rlabel metal1 -215 560 -215 560 1 Y
rlabel metal1 -215 646 -215 646 1 Y
rlabel metal2 -106 53 -106 53 1 X0
rlabel metal2 -114 53 -114 53 1 X1
rlabel metal2 -122 53 -122 53 1 X2
rlabel metal2 -130 53 -130 53 1 X3
rlabel metal2 -138 53 -138 53 1 X4
rlabel metal2 -146 53 -146 53 1 X5
rlabel metal2 -154 53 -154 53 1 X6
rlabel metal2 -162 53 -162 53 1 X7
<< end >>
