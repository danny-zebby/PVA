magic
tech scmos
timestamp 1715140968
<< metal1 >>
rect 996 2343 2605 2347
rect 2609 2343 2665 2347
rect 996 2335 2613 2339
rect 2617 2335 2665 2339
rect 996 2327 2621 2331
rect 2625 2327 2665 2331
rect 996 2319 2629 2323
rect 2633 2319 2665 2323
rect 996 2311 2637 2315
rect 2641 2311 2665 2315
rect 996 2303 2645 2307
rect 2649 2303 2665 2307
rect 996 2295 2653 2299
rect 2657 2295 2665 2299
rect 996 2287 2661 2291
rect 313 1911 351 1915
rect 321 1859 351 1863
rect 2541 1331 2571 1335
rect 2542 1279 2563 1283
rect 72 1113 101 1117
rect 1359 1026 1716 1030
rect 1720 1026 1721 1030
rect 1359 1018 1708 1022
rect 1712 1018 1721 1022
rect 1359 1010 1700 1014
rect 1704 1010 1721 1014
rect 1359 1002 1692 1006
rect 1696 1002 1721 1006
rect 1359 994 1684 998
rect 1688 994 1721 998
rect 1359 986 1676 990
rect 1680 986 1721 990
rect 1359 978 1668 982
rect 1672 978 1721 982
rect 1359 970 1660 974
rect 1664 970 1721 974
rect 2264 877 2571 881
rect 2238 825 2563 829
rect 10 36 14 40
rect 10 28 14 32
rect 10 20 14 24
rect 10 12 14 16
<< m2contact >>
rect 309 2592 313 2596
rect 317 2540 321 2544
rect 2605 2343 2609 2347
rect 2613 2335 2617 2339
rect 2621 2327 2625 2331
rect 2629 2319 2633 2323
rect 2637 2311 2641 2315
rect 2645 2303 2649 2307
rect 2653 2295 2657 2299
rect 2661 2287 2665 2291
rect 309 1911 313 1915
rect 317 1859 321 1863
rect 2571 1331 2575 1335
rect 2563 1279 2567 1283
rect 32 1136 36 1140
rect 1235 1123 1239 1127
rect 68 1113 72 1117
rect 101 1113 105 1117
rect 1227 1115 1231 1119
rect 1219 1107 1223 1111
rect 1211 1099 1215 1103
rect 1716 1026 1720 1030
rect 1708 1018 1712 1022
rect 1700 1010 1704 1014
rect 1692 1002 1696 1006
rect 1684 994 1688 998
rect 1676 986 1680 990
rect 1668 978 1672 982
rect 1660 970 1664 974
rect 2571 877 2575 881
rect 2563 825 2567 829
<< metal2 >>
rect 65 1615 69 2453
rect 101 1615 105 2496
rect 309 1915 313 2592
rect 317 1863 321 2540
rect 2605 2478 2609 2482
rect 2613 2478 2617 2482
rect 2621 2478 2625 2482
rect 2629 2478 2633 2482
rect 2637 2478 2641 2482
rect 2645 2478 2649 2482
rect 2653 2478 2657 2482
rect 2661 2478 2665 2482
rect 618 1185 622 1189
rect 32 868 36 1136
rect 101 1117 105 1179
rect 1211 1146 1215 1150
rect 273 1123 277 1127
rect 281 1123 285 1126
rect 289 1123 293 1126
rect 297 1122 301 1126
rect 68 868 72 1113
rect 1660 974 1664 1030
rect 1660 885 1664 970
rect 1668 982 1672 1030
rect 1668 885 1672 978
rect 1676 990 1680 1030
rect 1676 885 1680 986
rect 1684 998 1688 1030
rect 1684 885 1688 994
rect 1692 1006 1696 1030
rect 1692 885 1696 1002
rect 1700 1014 1704 1030
rect 1700 885 1704 1010
rect 1708 1022 1712 1030
rect 1708 885 1712 1018
rect 1716 885 1720 1026
rect 2563 829 2567 1279
rect 2571 881 2575 1331
rect 2605 1170 2609 2343
rect 2613 2339 2617 2347
rect 2613 1264 2617 2335
rect 2621 2331 2625 2347
rect 2621 1264 2625 2327
rect 2629 2323 2633 2347
rect 2629 1264 2633 2319
rect 2637 2315 2641 2347
rect 2637 1264 2641 2311
rect 2645 2307 2649 2347
rect 2645 1264 2649 2303
rect 2653 2299 2657 2347
rect 2653 1264 2657 2295
rect 2661 2291 2665 2347
rect 2661 1264 2665 2287
rect 2605 1161 2609 1165
rect 2613 1161 2617 1165
rect 2621 1161 2625 1165
rect 2629 1161 2633 1165
rect 2637 1161 2641 1165
rect 2645 1161 2649 1165
rect 2653 1161 2657 1165
rect 2661 1161 2665 1165
rect 2266 12 2270 16
rect 2274 12 2278 16
rect 2282 12 2286 16
rect 2290 12 2294 16
rect 2298 12 2302 16
rect 2306 12 2310 16
rect 2314 12 2318 16
rect 2322 12 2326 16
use VelocityDetector  VelocityDetector_0
timestamp 1715140639
transform 1 0 9 0 1 1156
box -20 -186 2656 1091
use VelocityDetector  VelocityDetector_1
timestamp 1715140639
transform 1 0 9 0 1 2473
box -20 -186 2656 1091
use pvaPosition  pvaPosition_0
timestamp 1715140639
transform 1 0 0 0 1 4
box 0 -4 2326 941
<< labels >>
rlabel metal1 12 30 12 30 1 RST
rlabel metal1 12 22 12 22 1 CLK
rlabel metal1 12 14 12 14 1 B
rlabel metal1 12 38 12 38 1 A
rlabel metal2 2655 1163 2655 1163 1 V1
rlabel metal2 2647 1163 2647 1163 1 V2
rlabel metal2 2639 1163 2639 1163 1 V3
rlabel metal2 2631 1163 2631 1163 1 V4
rlabel metal2 2663 1163 2663 1163 1 V0
rlabel metal2 2623 1163 2623 1163 1 V5
rlabel metal2 2615 1163 2615 1163 1 V6
rlabel metal2 2607 1163 2607 1163 1 V7
rlabel m2contact 2565 827 2565 827 1 VSS
rlabel m2contact 2573 879 2573 879 1 VDD
rlabel metal2 2324 14 2324 14 1 P7
rlabel metal2 2316 14 2316 14 1 P6
rlabel metal2 2308 14 2308 14 1 P5
rlabel metal2 2300 14 2300 14 1 P4
rlabel metal2 2292 14 2292 14 1 P3
rlabel metal2 2284 14 2284 14 1 P2
rlabel metal2 2276 14 2276 14 1 P1
rlabel metal2 2268 14 2268 14 1 P0
rlabel metal2 299 1124 299 1124 1 C0
rlabel metal2 291 1124 291 1124 1 C1
rlabel metal2 283 1124 283 1124 1 C2
rlabel metal2 275 1125 275 1125 1 C3
rlabel m2contact 1213 1101 1213 1101 1 X0
rlabel m2contact 1221 1109 1221 1109 1 X1
rlabel m2contact 1229 1117 1229 1117 1 X2
rlabel m2contact 1237 1125 1237 1125 1 X3
rlabel metal2 620 1187 620 1187 1 NOR4
rlabel metal2 2663 2480 2663 2480 7 A0
rlabel metal2 2655 2480 2655 2480 1 A1
rlabel metal2 2647 2480 2647 2480 1 A2
rlabel metal2 2639 2480 2639 2480 1 A3
rlabel metal2 2631 2480 2631 2480 1 A4
rlabel metal2 2623 2480 2623 2480 1 A5
rlabel metal2 2615 2480 2615 2480 1 A6
rlabel metal2 2607 2480 2607 2480 1 A7
<< end >>
