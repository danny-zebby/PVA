magic
tech scmos
timestamp 1712274593
<< nwell >>
rect -6 26 30 62
<< ntransistor >>
rect 7 8 9 12
rect 15 8 17 12
<< ptransistor >>
rect 7 32 9 48
rect 15 32 17 48
<< ndiffusion >>
rect 6 8 7 12
rect 9 8 10 12
rect 14 8 15 12
rect 17 8 18 12
<< pdiffusion >>
rect 6 32 7 48
rect 9 32 15 48
rect 17 32 18 48
<< ndcontact >>
rect 2 8 6 12
rect 10 8 14 12
rect 18 8 22 12
<< pdcontact >>
rect 2 32 6 48
rect 18 32 22 48
<< psubstratepcontact >>
rect 2 0 6 4
<< nsubstratencontact >>
rect 2 52 6 56
<< polysilicon >>
rect 7 48 9 50
rect 15 48 17 50
rect 7 20 9 32
rect 6 16 9 20
rect 7 12 9 16
rect 15 20 17 32
rect 15 16 18 20
rect 15 12 17 16
rect 7 6 9 8
rect 15 6 17 8
<< polycontact >>
rect 2 16 6 20
rect 18 16 22 20
<< metal1 >>
rect 0 52 2 56
rect 6 52 24 56
rect 2 48 6 52
rect 10 28 22 32
rect 10 12 14 28
rect 2 4 6 8
rect 18 4 22 8
rect 0 0 2 4
rect 6 0 24 4
<< labels >>
rlabel nsubstratencontact 4 54 4 54 1 VDD
rlabel polycontact 4 18 4 18 1 A
rlabel polycontact 20 18 20 18 1 B
rlabel psubstratepcontact 4 2 4 2 1 VSS
rlabel metal1 12 25 12 25 1 Y
<< end >>
