magic
tech scmos
timestamp 1711593098
<< nwell >>
rect 10 52 14 56
<< polycontact >>
rect 7 28 11 32
rect 27 28 31 32
rect 17 20 21 24
rect 37 20 41 24
<< metal1 >>
rect 10 52 14 56
rect 62 21 66 25
rect 46 16 54 20
rect 10 0 14 4
use INV  INV_0
timestamp 1711561836
transform 1 0 52 0 1 0
box -4 0 20 59
use NAND4  NAND4_0
timestamp 1711591893
transform 1 0 4 0 1 0
box -4 0 54 62
<< labels >>
rlabel metal1 64 23 64 23 1 Y
rlabel metal1 12 2 12 2 1 VSS
rlabel metal1 12 54 12 54 1 VDD
rlabel polycontact 9 30 9 30 1 A
rlabel polycontact 19 22 19 22 1 B
rlabel polycontact 29 30 29 30 1 C
rlabel polycontact 39 22 39 22 1 D
<< end >>
