magic
tech scmos
timestamp 1714413118
<< nwell >>
rect 117 58 129 62
<< metal1 >>
rect 0 52 6 56
rect 1 28 7 32
rect 0 20 17 24
rect 122 16 134 20
rect 162 15 166 21
rect 0 0 6 4
rect 0 -8 23 -4
rect 62 -10 146 -6
rect 0 -16 33 -12
rect 0 -24 67 -20
rect 0 -32 77 -28
rect 0 -40 87 -36
rect 0 -48 97 -44
<< m2contact >>
rect 23 24 27 28
rect 33 24 37 28
rect 67 24 71 28
rect 77 24 81 28
rect 87 24 91 28
rect 97 24 101 28
rect 146 20 150 24
rect 58 16 62 20
rect 23 -8 27 -4
rect 58 -10 62 -6
rect 146 -10 150 -6
rect 33 -16 37 -12
rect 67 -24 71 -20
rect 77 -32 81 -28
rect 87 -40 91 -36
rect 97 -48 101 -44
<< metal2 >>
rect 23 -4 27 24
rect 33 -12 37 24
rect 58 -6 62 16
rect 67 -20 71 24
rect 77 -28 81 24
rect 87 -36 91 24
rect 97 -44 101 24
rect 146 -6 150 20
use AND4  AND4_0
timestamp 1711593098
transform 1 0 -4 0 1 0
box 0 0 72 62
use AND4  AND4_1
timestamp 1711593098
transform 1 0 60 0 1 0
box 0 0 72 62
use OR2  OR2_0
timestamp 1712274593
transform 1 0 128 0 1 0
box -6 0 44 62
<< labels >>
rlabel metal1 1 54 1 54 3 VDD
rlabel metal1 2 30 2 30 1 A
rlabel metal1 1 22 1 22 3 B
rlabel metal1 1 2 1 2 3 VSS
rlabel metal1 1 -6 1 -6 3 C
rlabel metal1 1 -14 1 -14 3 D
rlabel metal1 1 -22 1 -22 3 E
rlabel metal1 1 -30 1 -30 3 F
rlabel metal1 1 -38 1 -38 3 G
rlabel metal1 1 -46 1 -46 2 H
rlabel metal1 164 18 164 18 1 Y
<< end >>
