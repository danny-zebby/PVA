magic
tech scmos
timestamp 1711564045
<< psubstratepcontact >>
rect 9 0 13 4
<< polycontact >>
rect 9 26 13 30
rect 19 26 23 30
<< metal1 >>
rect 12 52 16 56
rect 44 24 48 28
rect 29 16 36 20
use INV  INV_0
timestamp 1711561836
transform 1 0 34 0 1 0
box -4 0 20 59
use NAND2  NAND2_0
timestamp 1711563584
transform 1 0 6 0 1 0
box -6 0 34 62
<< labels >>
rlabel metal1 14 54 14 54 1 VDD
rlabel metal1 46 26 46 26 1 Y
rlabel polycontact 11 28 11 28 1 A
rlabel polycontact 21 28 21 28 1 B
rlabel psubstratepcontact 11 2 11 2 1 VSS
<< end >>
